`timescale 1ns/1ps
`default_nettype none

// ═══════════════════════════════════════════════════════════════════════════════
// PE Module Testbench - Professional Version
// Author: Chen Weidong
// Date: 2026-01-20
//
// Features:
// - FSDB waveform generation for Verdi
// - Self-checking test cases
// - Comprehensive test coverage
// - Clear pass/fail reporting
// ═══════════════════════════════════════════════════════════════════════════════

module tb_pe;

    // ═══════════════════════════════════════════════════════════════════════════
    // 信号声明
    // ═══════════════════════════════════════════════════════════════════════════

    logic clk;
    logic rst;

    // North wires (from above)
    logic signed [15:0] pe_psum_in;
    logic signed [15:0] pe_weight_in;
    logic pe_accept_w_in;

    // West wires (from left)
    logic signed [15:0] pe_input_in;
    logic pe_valid_in;
    logic pe_switch_in;
    logic pe_enabled;

    // South wires (to below)
    logic signed [15:0] pe_psum_out;
    logic signed [15:0] pe_weight_out;

    // East wires (to right)
    logic signed [15:0] pe_input_out;
    logic pe_valid_out;
    logic pe_switch_out;

    // 测试统计
    int test_count = 0;
    int pass_count = 0;
    int fail_count = 0;

    // 随机测试配置
    int random_test_num = 10;  // 随机测试数量

    // ═══════════════════════════════════════════════════════════════════════════
    // DUT 实例化
    // ═══════════════════════════════════════════════════════════════════════════

    pe #(
        .DATA_WIDTH(16)
    ) dut (
        .clk(clk),
        .rst(rst),
        .pe_psum_in(pe_psum_in),
        .pe_weight_in(pe_weight_in),
        .pe_accept_w_in(pe_accept_w_in),
        .pe_input_in(pe_input_in),
        .pe_valid_in(pe_valid_in),
        .pe_switch_in(pe_switch_in),
        .pe_enabled(pe_enabled),
        .pe_psum_out(pe_psum_out),
        .pe_weight_out(pe_weight_out),
        .pe_input_out(pe_input_out),
        .pe_valid_out(pe_valid_out),
        .pe_switch_out(pe_switch_out)
    );

    // ═══════════════════════════════════════════════════════════════════════════
    // 时钟生成 (10ns 周期 = 100MHz)
    // ═══════════════════════════════════════════════════════════════════════════

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // ═══════════════════════════════════════════════════════════════════════════
    // FSDB 波形生成（用于 Verdi 调试）
    // ═══════════════════════════════════════════════════════════════════════════

    initial begin
        // 从 build/ 目录到 waveforms/ 需要两层 ../
        // build/ -> ../ -> vcs/ -> ../ -> sim/ -> waveforms/
        $display("═══════════════════════════════════════════════════════════════════");
        $display("🔍 [DEBUG] 开始配置FSDB波形dump");
        $display("═══════════════════════════════════════════════════════════════════");

        $fsdbDumpfile("../../waveforms/tb_pe.fsdb");
        $display("✅ [DEBUG] fsdbDumpfile 已调用");

        // 官方推荐语法：depth=0表示dump所有层次
        $fsdbDumpvars(0, tb_pe);
        $display("✅ [DEBUG] fsdbDumpvars(0, tb_pe) 已调用");
        $display("═══════════════════════════════════════════════════════════════════\n");
    end

    // ═══════════════════════════════════════════════════════════════════════════
    // 断言（Assertion）- 为 UVM 验证做准备
    // ═══════════════════════════════════════════════════════════════════════════

    // 断言1：复位期间输出应该为0
    // 注意：复位是同步复位，需要在复位后的下一个时钟周期检查
    property reset_output_zero;
        @(posedge clk) (rst) |=> (pe_psum_out == 0);
    endproperty
    assert property (reset_output_zero)
        else $error("[ASSERTION FAIL] 复位后输出不为0!");

    // 断言2：数据传播检查 - valid信号传播到输出
    // 注意：在脉动阵列中，valid可以连续多周期保持高电平，这是正常的
    property valid_propagation;
        @(posedge clk) disable iff (rst)
            pe_valid_in |-> ##1 pe_valid_out;
    endproperty
    assert property (valid_propagation)
        else $warning("[ASSERTION WARN] valid 信号未正确传播到输出!");

    // ═══════════════════════════════════════════════════════════════════════════
    // Q8.8 定点数转换函数
    // ═══════════════════════════════════════════════════════════════════════════

    function automatic logic [15:0] to_fixed(real val);
        return $signed($rtoi(val * 256.0)) & 16'hFFFF;
    endfunction

    function automatic real from_fixed(logic [15:0] val);
        logic signed [15:0] signed_val;
        signed_val = val;
        return $itor(signed_val) / 256.0;
    endfunction

    // ═══════════════════════════════════════════════════════════════════════════
    // 测试任务
    // ═══════════════════════════════════════════════════════════════════════════

    task automatic reset_dut();
        $display("[%0t] 🔄 复位 DUT", $time);
        rst = 1;
        pe_enabled = 0;
        pe_valid_in = 0;
        pe_accept_w_in = 0;
        pe_switch_in = 0;
        pe_input_in = 16'h0000;
        pe_weight_in = 16'h0000;
        pe_psum_in = 16'h0000;

        repeat(3) @(posedge clk);
        rst = 0;
        pe_enabled = 1;
        @(posedge clk);
        $display("[%0t] ✅ 复位完成\n", $time);
    endtask

    task automatic load_weight(real weight_val);
        $display("[%0t] 📥 加载权重: %.2f", $time, weight_val);
        pe_accept_w_in = 1;
        pe_weight_in = to_fixed(weight_val);
        @(posedge clk);
        pe_accept_w_in = 0;
        $display("[%0t] ✅ 权重已加载到后台寄存器", $time);
    endtask

    task automatic switch_weight();
        $display("[%0t] 🔄 切换权重（后台→前台）", $time);
        pe_switch_in = 1;
        @(posedge clk);
        pe_switch_in = 0;
        @(posedge clk);  // 等待切换完成（纯时序逻辑需要1周期）
        $display("[%0t] ✅ 权重切换完成", $time);
    endtask

    task automatic mac_operation(
        input real input_val,
        input real psum_val,
        input real expected_out,
        input string test_name
    );
        real actual_out;
        real error;

        test_count++;
        $display("[%0t] 🧮 MAC 运算 [%s]: %.2f * weight + %.2f",
                 $time, test_name, input_val, psum_val);

        // 设置输入数据和valid信号
        pe_input_in = to_fixed(input_val);
        pe_psum_in = to_fixed(psum_val);
        pe_valid_in = 1;

        // 工业级验证标准做法：等待2个时钟周期
        // T1: PE捕获输入数据
        @(posedge clk);

        // T2: PE输出计算结果（流水线延迟）
        @(posedge clk);

        // 在T2时钟沿之后采样，此时输出已经稳定
        actual_out = from_fixed(pe_psum_out);
        error = $abs(actual_out - expected_out);

        // 采样完成后拉低valid信号
        pe_valid_in = 0;

        $display("[%0t] 📊 期望: %.4f, 实际: %.4f, 误差: %.4f (0x%04h)",
                 $time, expected_out, actual_out, error, pe_psum_out);

        // Q8.8 定点数精度约为 1/256 ≈ 0.0039
        // 考虑到乘法累积误差，设置容差为 0.02（约5个LSB）
        if (error < 0.02) begin
            $display("[%0t] ✅ PASS\n", $time);
            pass_count++;
        end else begin
            $display("[%0t] ❌ FAIL - 误差超出容差范围!\n", $time);
            fail_count++;
        end
    endtask

    // ═══════════════════════════════════════════════════════════════════════════
    // 随机测试任务（为 UVM 做准备）
    // ═══════════════════════════════════════════════════════════════════════════
    task automatic random_mac_test(input int num_tests, input real weight_val);
        real rand_input, rand_psum, expected;
        int seed = $urandom();  // 随机种子

        $display("[%0t] 🎲 开始随机测试 (%0d 次)", $time, num_tests);
        $display("[%0t] 🔑 随机种子: %0d", $time, seed);

        load_weight(weight_val);
        switch_weight();

        for (int i = 0; i < num_tests; i++) begin
            // 生成随机数（范围：-2.0 ~ 2.0）
            // 限制范围以避免超出 Q8.8 表示范围（-128 ~ 127.996）
            // 对于 weight=1.5，最大输出约为 2.0*1.5+2.0=5.0，安全范围内
            rand_input = ($urandom_range(0, 400) - 200) / 100.0;
            rand_psum = ($urandom_range(0, 400) - 200) / 100.0;

            // 计算期望值
            expected = rand_input * weight_val + rand_psum;

            // 检查是否超出 Q8.8 表示范围
            if (expected > 127.0 || expected < -128.0) begin
                $display("[%0t] ⚠️  跳过测试-%0d: 期望值 %.4f 超出 Q8.8 范围",
                         $time, i+1, expected);
                continue;
            end

            // 执行 MAC 运算
            mac_operation(rand_input, rand_psum, expected,
                         $sformatf("随机测试-%0d", i+1));
        end

        $display("[%0t] ✅ 随机测试完成\n", $time);
    endtask

    // ═══════════════════════════════════════════════════════════════════════════
    // 主测试流程
    // ═══════════════════════════════════════════════════════════════════════════

    initial begin
        $display("═══════════════════════════════════════════════════════════════════");
        $display("🧪 PE Module Testbench - Professional Version");
        $display("═══════════════════════════════════════════════════════════════════");
        $display("测试内容:");
        $display("  1. 权重加载到后台寄存器");
        $display("  2. 权重切换到前台寄存器");
        $display("  3. MAC 运算验证 (5个定向测试)");
        $display("  4. 随机测试 (%0d 次)", random_test_num);
        $display("  5. 断言检查（Assertion）");
        $display("═══════════════════════════════════════════════════════════════════\n");

        // ═══════════════════════════════════════════════════════════════════════
        // Test 1: 基础 MAC 运算
        // ═══════════════════════════════════════════════════════════════════════
        $display("[Test 1] 基础 MAC 运算");
        $display("───────────────────────────────────────────────────────────────────");

        reset_dut();
        load_weight(2.0);
        switch_weight();
        mac_operation(3.0, 1.0, 7.0, "基础运算");

        // ═══════════════════════════════════════════════════════════════════════
        // Test 2: 零值测试
        // ═══════════════════════════════════════════════════════════════════════
        $display("[Test 2] 零值测试");
        $display("───────────────────────────────────────────────────────────────────");

        reset_dut();
        load_weight(0.0);
        switch_weight();
        mac_operation(5.0, 0.0, 0.0, "零权重");

        // ═══════════════════════════════════════════════════════════════════════
        // Test 3: 负数测试
        // ═══════════════════════════════════════════════════════════════════════
        $display("[Test 3] 负数测试");
        $display("───────────────────────────────────────────────────────────────────");

        reset_dut();
        load_weight(-1.5);
        switch_weight();
        mac_operation(2.0, 4.0, 1.0, "负权重");

        // ═══════════════════════════════════════════════════════════════════════
        // Test 4: 小数精度测试
        // ═══════════════════════════════════════════════════════════════════════
        $display("[Test 4] 小数精度测试");
        $display("───────────────────────────────────────────────────────────────────");

        reset_dut();
        load_weight(0.5);
        switch_weight();
        mac_operation(1.25, 0.25, 0.875, "小数精度");

        // ═══════════════════════════════════════════════════════════════════════
        // Test 5: 连续 MAC 运算
        // ═══════════════════════════════════════════════════════════════════════
        $display("[Test 6] 连续 MAC 运算");
        $display("───────────────────────────────────────────────────────────────────");

        reset_dut();
        load_weight(1.0);
        switch_weight();
        mac_operation(1.0, 0.0, 1.0, "连续-1");
        mac_operation(2.0, 0.0, 2.0, "连续-2");
        mac_operation(3.0, 0.0, 3.0, "连续-3");

        // ═══════════════════════════════════════════════════════════════════════
        // Test 6: 随机测试（新增！）
        // ═══════════════════════════════════════════════════════════════════════
        $display("[Test 6] 随机测试");
        $display("───────────────────────────────────────────────────────────────────");

        reset_dut();
        random_mac_test(random_test_num, 1.5);  // 权重=1.5，运行10次随机测试

        // ═══════════════════════════════════════════════════════════════════════
        // 测试完成 - 打印统计信息
        // ═══════════════════════════════════════════════════════════════════════

        repeat(10) @(posedge clk);

        $display("═══════════════════════════════════════════════════════════════════");
        $display("📊 测试统计");
        $display("═══════════════════════════════════════════════════════════════════");
        $display("  总测试数: %0d", test_count);
        $display("  通过数:   %0d", pass_count);
        $display("  失败数:   %0d", fail_count);
        $display("  通过率:   %.1f%%", (pass_count * 100.0) / test_count);
        $display("═══════════════════════════════════════════════════════════════════");

        if (fail_count == 0) begin
            $display("✅ 所有测试通过!");
            $display("═══════════════════════════════════════════════════════════════════\n");
            $finish(0);  // 返回 0 表示成功
        end else begin
            $display("❌ 有 %0d 个测试失败!", fail_count);
            $display("═══════════════════════════════════════════════════════════════════\n");
            $finish(1);  // 返回 1 表示失败
        end
    end

    // ═══════════════════════════════════════════════════════════════════════════
    // 超时保护
    // ═══════════════════════════════════════════════════════════════════════════

    initial begin
        #10000;  // 10us 超时
        $display("\n❌ 测试超时!");
        $display("═══════════════════════════════════════════════════════════════════\n");
        $finish(2);  // 返回 2 表示超时
    end

endmodule

`default_nettype wire
